// Code for nand gate
module nand_gate(
  input a,
  input b,
  output y
);
 nand(y,a,b);
 endmodule
